module app ( 
    output wire led
); 
 
assign led = 1'b1; 

endmodule 
